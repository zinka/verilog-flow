// This is a simple example.
// 
// 
//
//		
//
// -----------------------------------------------------------------------------
// Copyright (c) 2014-2020 All rights reserved
// -----------------------------------------------------------------------------
// Author : Srinivasa Rao Zinka (zinka) srinivas.zinka@gmail.com
// File   : top.v
// Create : 2020-04-23 08:27:08
// Revise : 2020-04-23 11:00:32
// Editor : sublime text3, tab size (4)
// -----------------------------------------------------------------------------


// `define ENABLE_ADC_CLOCK
// `define ENABLE_CLOCK1
// `define ENABLE_CLOCK2
// `define ENABLE_SDRAM
// `define ENABLE_HEX0
// `define ENABLE_HEX1
// `define ENABLE_HEX2
// `define ENABLE_HEX3
// `define ENABLE_HEX4
// `define ENABLE_HEX5
// `define ENABLE_KEY
// `define ENABLE_LED
// `define ENABLE_SW
// `define ENABLE_VGA
// `define ENABLE_ACCELEROMETER
// `define ENABLE_ARDUINO
// `define ENABLE_GPIO

module top (
	//////////// ADC CLOCK: 3.3-V LVTTL //////////
	`ifdef ENABLE_ADC_CLOCK
	input         ADC_CLK_10     ,
	`endif
	//////////// CLOCK 1: 3.3-V LVTTL //////////
	`ifdef ENABLE_CLOCK1
	input         MAX10_CLK1_50  ,
	`endif
	//////////// CLOCK 2: 3.3-V LVTTL //////////
	`ifdef ENABLE_CLOCK2
	input         MAX10_CLK2_50  ,
	`endif
	//////////// SDRAM: 3.3-V LVTTL //////////
	`ifdef ENABLE_SDRAM
	output [12:0] DRAM_ADDR      ,
	output [ 1:0] DRAM_BA        ,
	output        DRAM_CAS_N     ,
	output        DRAM_CKE       ,
	output        DRAM_CLK       ,
	output        DRAM_CS_N      ,
	inout  [15:0] DRAM_DQ        ,
	output        DRAM_LDQM      ,
	output        DRAM_RAS_N     ,
	output        DRAM_UDQM      ,
	output        DRAM_WE_N      ,
	`endif
	//////////// SEG7: 3.3-V LVTTL //////////
	`ifdef ENABLE_HEX0
	output [ 7:0] HEX0           ,
	`endif
	`ifdef ENABLE_HEX1
	output [ 7:0] HEX1           ,
	`endif
	`ifdef ENABLE_HEX2
	output [ 7:0] HEX2           ,
	`endif
	`ifdef ENABLE_HEX3
	output [ 7:0] HEX3           ,
	`endif
	`ifdef ENABLE_HEX4
	output [ 7:0] HEX4           ,
	`endif
	`ifdef ENABLE_HEX5
	output [ 7:0] HEX5           ,
	`endif
	//////////// KEY: 3.3 V SCHMITT TRIGGER //////////
	`ifdef ENABLE_KEY
	input  [ 1:0] KEY            ,
	`endif
	//////////// LED: 3.3-V LVTTL //////////
	`ifdef ENABLE_LED
	output [ 9:0] LEDR           ,
	`endif
	//////////// SW: 3.3-V LVTTL //////////
	`ifdef ENABLE_SW
	input  [ 9:0] SW             ,
	`endif
	//////////// VGA: 3.3-V LVTTL //////////
	`ifdef ENABLE_VGA
	output [ 3:0] VGA_B          ,
	output [ 3:0] VGA_G          ,
	output        VGA_HS         ,
	output [ 3:0] VGA_R          ,
	output        VGA_VS         ,
	`endif
	//////////// Accelerometer: 3.3-V LVTTL //////////
	`ifdef ENABLE_ACCELEROMETER
	output        GSENSOR_CS_N   ,
	input  [ 2:1] GSENSOR_INT    ,
	output        GSENSOR_SCLK   ,
	inout         GSENSOR_SDI    ,
	inout         GSENSOR_SDO    ,
	`endif
	//////////// Arduino: 3.3-V LVTTL //////////
	`ifdef ENABLE_ARDUINO
	inout  [15:0] ARDUINO_IO     ,
	inout         ARDUINO_RESET_N,
	`endif
	//////////// GPIO, GPIO connect to GPIO Default: 3.3-V LVTTL //////////
	`ifdef ENABLE_GPIO
	inout  [35:0] GPIO
	`endif
);





endmodule
